** Profile: "SCHEMATIC1-SeniorDesign2"  [ U:\SeniorDesign\Orcad\seniordesign2-pspicefiles\schematic1\seniordesign2.sim ] 

** Creating circuit file "SeniorDesign2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "U:\SeniorDesign\Orcad\sboma53\OPA4830.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 
.OPTIONS ADVCONV
.OPTIONS VNTOL= 100n
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
